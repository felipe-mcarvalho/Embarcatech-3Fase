module aes_round (
    input  wire [127:0] state_in,      // Dados de entrada da rodada
    input  wire [127:0] round_key,     // A chave espec�fica desta rodada
    input  wire         is_last_round, // 0 = Rodada Normal, 1 = �ltima rodada 
    output wire [127:0] state_out      // Dados de sa�da
);

    // Fios internos para conectar os blocos
    wire [127:0] after_subbytes;
    wire [127:0] after_shiftrows;
    wire [127:0] after_mixcolumns;
    
    // Inst�ncia subBytes
    aes_sub_bytes u_subbytes (
        .state_in  (state_in),
        .state_out (after_subbytes)
    );

    // Inst�ncia shiftRows
    aes_shift_rows u_shiftrows (
        .state_in  (after_subbytes),
        .state_out (after_shiftrows)
    );

    // Inst�ncia mixColumns
    aes_mix_columns u_mixcolumns (
        .state_in  (after_shiftrows),
        .state_out (after_mixcolumns)
    );


    // L�gica do MUX para a �ltima rodada
    // Se for a �ltima rodada, pegar o dado  do ShiftRows.
    // Se for rodada normal,   pegar o dado do MixColumns.
	    
    wire [127:0] mix_mux_out; // Fio que decide quem entra no AddRoundKey
    assign mix_mux_out = (is_last_round) ? after_shiftrows : after_mixcolumns;


    // Inst�ncia addRoundKey
    aes_add_round_key u_addroundkey (
        .state_in  (mix_mux_out),
        .round_key (round_key),
        .state_out (state_out)
    );

endmodule